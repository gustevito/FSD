--------------------------------------
-- Biblioteca
--------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

--------------------------------------
-- Entidade
--------------------------------------
entity desafio is
    port( --COMPLETAR
        );
end entity;

--------------------------------------
-- Arquitetura
--------------------------------------
architecture behaviour of desafio is
  --COMPLETAR
begin                           
  
  --COMPLETAR

end architecture;