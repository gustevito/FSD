--------------------------------------
-- Biblioteca
--------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;

--------------------------------------
-- Entidade
--------------------------------------
entity ex3 is
  port( -- <COMPLETAR>
      );
end entity;

--------------------------------------
-- Arquitetura
--------------------------------------
architecture ex3 of ex3 is
  -- <COMPLETAR>
begin

  sd <= -- <COMPLETAR>
	
  BB <= -- <COMPLETAR>
	
end architecture;