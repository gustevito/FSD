--------------------------------------
-- Biblioteca
--------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;

--------------------------------------
-- Entidade
--------------------------------------
entity ex2 is
  port( -- <COMPLETAR>
      );
end entity;

--------------------------------------
-- Arquitetura
--------------------------------------
architecture ex2 of ex2 is
begin
  -- <COMPLETAR>
end architecture;