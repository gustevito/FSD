--------------------------------------
-- Biblioteca
--------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

--------------------------------------
-- Entidade
--------------------------------------
entity ex1 is        
    port( -- <COMPLETAR>
        );
end entity;

--------------------------------------
-- Arquitetura
--------------------------------------
architecture ex1 of ex1 is    
    -- <COMPLETAR>
begin 

    -- <COMPLETAR>

end architecture;