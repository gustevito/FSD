--------------------------------------
-- Biblioteca
--------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

--------------------------------------
-- Entidade
--------------------------------------
entity ex_prova is        
    port( -- <COMPLETAR>
        );
end entity;

--------------------------------------
-- Arquitetura
--------------------------------------
architecture ex_prova of ex_prova is    
    -- <COMPLETAR>
begin 

    -- <COMPLETAR>

end architecture;