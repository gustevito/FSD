--------------------------------------
-- Biblioteca
--------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

--------------------------------------
-- Entidade
--------------------------------------
entity ex2 is        
    port( -- <COMPLETAR>
        );
end entity;

--------------------------------------
-- Arquitetura
--------------------------------------
architecture ex2 of ex2 is    
    -- <COMPLETAR>
begin 

    -- <COMPLETAR>

end architecture;