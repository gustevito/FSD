--------------------------------------
-- Biblioteca
--------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

--------------------------------------
-- Entidade
--------------------------------------
entity exercicio_avancado is        
    port( --COMPLETAR--
         );
end entity;

--------------------------------------
-- Arquitetura
--------------------------------------
architecture behavioral of exercicio_avancado is    
    --COMPLETAR--
begin 

    --COMPLETAR--

end architecture;