--------------------------------------
-- Biblioteca
--------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

--------------------------------------
-- Entidade
--------------------------------------
entity ex3 is        
    port( -- <COMPLETAR>
        );
end entity;

--------------------------------------
-- Arquitetura
--------------------------------------
architecture ex3 of ex3 is    
    -- <COMPLETAR>
begin 

    -- <COMPLETAR>

end architecture;